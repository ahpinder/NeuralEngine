package core_pkg;
    typedef enum af_control [3:0] {   //Signal to Control the activation Function
        ReLu = 4'b0000,
    }
endpackage